// File name:   key_expansion.sv
// Created:     4/19/2018
// Author:      Ryan Devlin
// Lab Section: 337-05
// Version:     1.0  Initial Design Entry
// Description: Turns a 128-bit key into a 1408-bit key.
`timescale 1ns / 100ps

module key_expansion
(
	input logic clk,
	input logic n_rst,
	input logic start_key_exp,
	input logic [127:0] key,
	output logic key_expanded,
	output logic [1407:0] exp_key
);

typedef enum bit [3:0] {IDLE, STATE_0, STATE_1, STATE_2, STATE_3, STATE_4, STATE_5, STATE_6, STATE_7, STATE_8, STATE_9, STATE_10} stateType;
stateType state, next_state;

logic [127:0] next_curr_key, curr_key;
logic [127:0] next_prev_key, prev_key;
logic [1407:0] next_exp_key;

logic [3:0] round_number;
logic [31:0] core_out;

keyScheduleCore U1 
(
	.inputWord(prev_key[31:0]), 
	.roundNumber(round_number), 
	.outputWord(core_out)
);

always_comb begin 
	next_state = state;

	case(state)
	IDLE: begin
		if(start_key_exp == 1'b1) begin
			next_state = STATE_0;
		end	
	end
	STATE_0: begin
		next_state = STATE_1;
	end
	STATE_1: begin
		next_state = STATE_2;
	end
	STATE_2: begin
		next_state = STATE_3;
	end
	STATE_3: begin
		next_state = STATE_4;
	end
	STATE_4: begin
		next_state = STATE_5;
	end
	STATE_5: begin
		next_state = STATE_6;
	end
	STATE_6: begin
		next_state = STATE_7;
	end
	STATE_7: begin
		next_state = STATE_8;
	end
	STATE_8: begin
		next_state = STATE_9;
	end
	STATE_9: begin
		next_state = STATE_10;
	end
	STATE_10: begin
		next_state = IDLE;
	end
	endcase
end

always_comb begin 
	next_curr_key = curr_key;
	next_prev_key = prev_key;
	next_exp_key = exp_key;
	key_expanded = 1'b0;
	round_number = 4'h0;	

	case(state)
	IDLE: begin
		next_curr_key = curr_key;
		next_prev_key = prev_key;
		next_exp_key = exp_key;
	end
	STATE_0: begin
		next_curr_key = curr_key;
		next_prev_key = key;
		next_exp_key[1407:1280] = key;
		round_number = 4'h0;
	end
	STATE_1: begin
		next_curr_key[127:96] = prev_key[127:96] ^ core_out;
		next_curr_key[95:64] = prev_key[95:64] ^ next_curr_key[127:96];
		next_curr_key[63:32] = prev_key[63:32] ^ next_curr_key[95:64];
		next_curr_key[31:0] = prev_key[31:0] ^ next_curr_key[63:32];
		next_prev_key = next_curr_key;
		next_exp_key[1279:1152] = next_curr_key;
		round_number = 4'h0;
	end
	STATE_2: begin
		next_curr_key[127:96] = prev_key[127:96] ^ core_out;
		next_curr_key[95:64] = prev_key[95:64] ^ next_curr_key[127:96];
		next_curr_key[63:32] = prev_key[63:32] ^ next_curr_key[95:64];
		next_curr_key[31:0] = prev_key[31:0] ^ next_curr_key[63:32];
		next_prev_key = next_curr_key;
		next_exp_key[1151:1024] = next_curr_key;
		round_number = 4'h1;
	end
	STATE_3: begin
		next_curr_key[127:96] = prev_key[127:96] ^ core_out;
		next_curr_key[95:64] = prev_key[95:64] ^ next_curr_key[127:96];
		next_curr_key[63:32] = prev_key[63:32] ^ next_curr_key[95:64];
		next_curr_key[31:0] = prev_key[31:0] ^ next_curr_key[63:32];
		next_prev_key = next_curr_key;
		next_exp_key[1023:896] = next_curr_key;
		round_number = 4'h2;
	end
	STATE_4: begin
		next_curr_key[127:96] = prev_key[127:96] ^ core_out;
		next_curr_key[95:64] = prev_key[95:64] ^ next_curr_key[127:96];
		next_curr_key[63:32] = prev_key[63:32] ^ next_curr_key[95:64];
		next_curr_key[31:0] = prev_key[31:0] ^ next_curr_key[63:32];
		next_prev_key = next_curr_key;
		next_exp_key[895:768] = next_curr_key;
		round_number = 4'h3;
	end
	STATE_5: begin
		next_curr_key[127:96] = prev_key[127:96] ^ core_out;
		next_curr_key[95:64] = prev_key[95:64] ^ next_curr_key[127:96];
		next_curr_key[63:32] = prev_key[63:32] ^ next_curr_key[95:64];
		next_curr_key[31:0] = prev_key[31:0] ^ next_curr_key[63:32];
		next_prev_key = next_curr_key;
		next_exp_key[767:640] = next_curr_key;
		round_number = 4'h4;
	end
	STATE_6: begin
		next_curr_key[127:96] = prev_key[127:96] ^ core_out;
		next_curr_key[95:64] = prev_key[95:64] ^ next_curr_key[127:96];
		next_curr_key[63:32] = prev_key[63:32] ^ next_curr_key[95:64];
		next_curr_key[31:0] = prev_key[31:0] ^ next_curr_key[63:32];
		next_prev_key = next_curr_key;
		next_exp_key[639:512] = next_curr_key;
		round_number = 4'h5;
	end
	STATE_7: begin
		next_curr_key[127:96] = prev_key[127:96] ^ core_out;
		next_curr_key[95:64] = prev_key[95:64] ^ next_curr_key[127:96];
		next_curr_key[63:32] = prev_key[63:32] ^ next_curr_key[95:64];
		next_curr_key[31:0] = prev_key[31:0] ^ next_curr_key[63:32];
		next_prev_key = next_curr_key;
		next_exp_key[511:384] = next_curr_key;
		round_number = 4'h6;
	end
	STATE_8: begin
		next_curr_key[127:96] = prev_key[127:96] ^ core_out;
		next_curr_key[95:64] = prev_key[95:64] ^ next_curr_key[127:96];
		next_curr_key[63:32] = prev_key[63:32] ^ next_curr_key[95:64];
		next_curr_key[31:0] = prev_key[31:0] ^ next_curr_key[63:32];
		next_prev_key = next_curr_key;
		next_exp_key[383:256] = next_curr_key;
		round_number = 4'h7;
	end
	STATE_9: begin
		next_curr_key[127:96] = prev_key[127:96] ^ core_out;
		next_curr_key[95:64] = prev_key[95:64] ^ next_curr_key[127:96];
		next_curr_key[63:32] = prev_key[63:32] ^ next_curr_key[95:64];
		next_curr_key[31:0] = prev_key[31:0] ^ next_curr_key[63:32];
		next_prev_key = next_curr_key;
		next_exp_key[255:128] = next_curr_key;
		round_number = 4'h8;
	end
	STATE_10: begin
		next_curr_key[127:96] = prev_key[127:96] ^ core_out;
		next_curr_key[95:64] = prev_key[95:64] ^ next_curr_key[127:96];
		next_curr_key[63:32] = prev_key[63:32] ^ next_curr_key[95:64];
		next_curr_key[31:0] = prev_key[31:0] ^ next_curr_key[63:32];
		next_prev_key = next_curr_key;
		next_exp_key[127:0] = next_curr_key;
		round_number = 4'h9;
		key_expanded = 1'b1;
	end
	endcase
end

always_ff @ (posedge clk, negedge n_rst) begin
	if(n_rst == 0) begin
		curr_key <= '0;
		prev_key <= '0;
		exp_key <= '0;
		state <= IDLE;
	end
	else begin
		curr_key <= next_curr_key;
		prev_key <= next_prev_key;
		exp_key <= next_exp_key;
		state <= next_state;
	end
end

endmodule
